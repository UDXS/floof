/*
Anf Floof
32-bit Embedded 3D Graphics Processor

Texture Color Parser
*/

module anfFl_tex_parser
	(
		input			reset,
		input			clk,
	);